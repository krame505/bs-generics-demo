
import "BDPI" function ActionValue#(Int#(32)) rxClient();
import "BDPI" function Action txClient(Bit#(8) data);
import "BDPI" function ActionValue#(Int#(32)) rxSim();
import "BDPI" function Action txSim(Bit#(8) data);
