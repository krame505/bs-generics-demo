-- Copyright 2021 Google LLC
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--      http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.

package UARTDemo where

import UART
import GetPut

interface UARTDemo =
  tx :: Bit 1 {-# always_ready, always_enabled #-}
  rx :: Bit 1 -> Action {-# always_ready, always_enabled, prefix="", arg_names = [rx] #-}

{-# verilog mkUARTDemo #-}
mkUARTDemo :: Module UARTDemo
mkUARTDemo = module
  uart <- mkUART 9600

  rules
    "echo": when True ==> do
       c <- uart.rxData.get
       uart.txData.put $ c + 1

  interface
    tx = uart.tx
    rx = uart.rx
