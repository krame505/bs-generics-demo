-- Copyright 2021 Google LLC
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--      http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.

package Counter where

import CShow
import Vector
import FIFO
import GetPut

type Id = Bit 16 -- Try changing the size

-- Try adding/reordering constructors
data CounterCommand = Num { id :: Id; val :: Int 32; }
                    | ResetSum (Int 32)
                    | ResetSquareSum (Int 64)
  deriving (Bits)

struct Result a =
  id :: Id
  val :: a
 deriving (Bits)

interface Counter =
  command :: Put CounterCommand
  sum :: Get (Result (Int 32))
  squareSum :: Get (Result (Int 64))

{-# verilog mkCounter #-}
mkCounter :: Module Counter
mkCounter = module
  commands <- mkFIFO
  sums <- mkFIFO
  squareSums <- mkFIFO

  sum :: Reg (Int 32) <- mkReg 0
  squareSum :: Reg (Int 64) <- mkReg 1

  rules
    "handle_command": when True ==> do
      -- $display "Handling command " (cshow c)
      case commands.first of
        Num { id = id; val = val; } -> do
          let newSum = sum + val
          let newSquareSum = squareSum + (signExtend val) * (signExtend val)
          sums.enq (Result { id = id; val = newSum; })
          squareSums.enq (Result { id = id; val = newSquareSum; })
          sum := newSum
          squareSum := newSquareSum
        ResetSum val -> do
          sum := val
        ResetSquareSum val -> do
          squareSum := val
      commands.deq

  interface
    command = toPut commands
    sum = toGet sums
    squareSum = toGet squareSums
