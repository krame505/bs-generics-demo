package UARTDemo where

import UART
import GetPut

interface UARTDemo =
  tx :: Bit 1 {-# always_ready, always_enabled #-}

{-# verilog mkUARTDemo #-}
mkUARTDemo :: Module UARTDemo
mkUARTDemo = module
  uart <- mkUART 9600

  i :: Reg (UInt 8) <- mkReg 0
  rules
    "put_demo": when True ==> do
       i := (i + 1) % 26
       uart.txData.put $ pack $ i + 65

  interface
    tx = uart.tx
