package Counter where

import CShow
import Vector
import FIFO
import GetPut

type Id = Bit 16 -- Try changing the size

-- Try adding/reordering constructors
data Command = Num { id :: Id; val :: Int 16; }
             | ResetSum (Int 16)
             | ResetProduct (Int 64)
  deriving (Bits)

struct Result a =
  id :: Id
  val :: a
 deriving (Bits)

interface Counter =
  command :: Put Command
  sum :: Get (Result (Int 16))
  product :: Get (Result (Int 64))

{-# verilog mkCounter #-}
mkCounter :: Module Counter
mkCounter = module
  commands <- mkFIFO
  sums <- mkFIFO
  products <- mkFIFO

  sum :: Reg (Int 16) <- mkReg 0
  product :: Reg (Int 64) <- mkReg 1

  rules
    "handle_command": when True ==> do
      -- $display "Handling command " (cshow c)
      case commands.first of
        Num { id = id; val = val; } -> do
          let newSum = sum + val
          let newProduct = product * signExtend val
          sums.enq (Result { id = id; val = newSum; })
          products.enq (Result { id = id; val = newProduct; })
          sum := newSum
          product := newProduct
        ResetSum val -> do
          sum := val
        ResetProduct val -> do
          product := val
      commands.deq

  interface
    command = toPut commands
    sum = toGet sums
    product = toGet products
