package Counter where

import CShow
import Vector
import FIFO
import GetPut

type Id = Bit 16 -- Try changing the size

-- Try adding/reordering constructors
data CounterCommand = Num { id :: Id; val :: Int 16; }
                    | ResetSum (Int 16)
                    | ResetSquareSum (Int 64)
  deriving (Bits)

struct Result a =
  id :: Id
  val :: a
 deriving (Bits)

interface Counter =
  command :: Put CounterCommand
  sum :: Get (Result (Int 16))
  squareSum :: Get (Result (Int 64))

{-# verilog mkCounter #-}
mkCounter :: Module Counter
mkCounter = module
  commands <- mkFIFO
  sums <- mkFIFO
  squareSums <- mkFIFO

  sum :: Reg (Int 16) <- mkReg 0
  squareSum :: Reg (Int 64) <- mkReg 1

  rules
    "handle_command": when True ==> do
      -- $display "Handling command " (cshow c)
      case commands.first of
        Num { id = id; val = val; } -> do
          let newSum = sum + val
          let newSquareSum = squareSum + (signExtend val) * (signExtend val)
          sums.enq (Result { id = id; val = newSum; })
          squareSums.enq (Result { id = id; val = newSquareSum; })
          sum := newSum
          squareSum := newSquareSum
        ResetSum val -> do
          sum := val
        ResetSquareSum val -> do
          squareSum := val
      commands.deq

  interface
    command = toPut commands
    sum = toGet sums
    squareSum = toGet squareSums
