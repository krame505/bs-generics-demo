package DemoSim where

import DemoSimIface
import Demo
import UART
import RGB
import Buttons

import GetPut
import Connectable
import FIFO

{-# verilog sysDemoSim #-}
sysDemoSim :: Module Empty
sysDemoSim = module
  demo <- mkDemo

  init <- mkReg False

  rules
    "tx": when True ==> do
      c <- demo.txData.get
      $display "Tx %x" c
      txData c

    "rx": when True ==> do
      c <- rxData
      if c /= negate 1
        then do $display "Rx %x" c
                demo.rxData.put $ truncate $ pack c
        else noAction
