package RGB where

import GetPut

struct RGB =
  red :: UInt 8
  green :: UInt 8
  blue :: UInt 8
 deriving (Bits)

interface RGBControl =
  state :: Put RGB
  red :: Bit 1 {-# always_ready, always_enabled #-}
  green :: Bit 1 {-# always_ready, always_enabled #-}
  blue :: Bit 1 {-# always_ready, always_enabled #-}

{-# verilog mkRGBControl #-}
mkRGBControl :: Module RGBControl
mkRGBControl = module
  state :: Reg RGB <- mkReg $ RGB {red = 0; green = 0; blue = 0;}
  count :: Reg (UInt 8) <- mkReg 0

  rules
    "update_count": when True ==> count := count + 1

  interface
    state = toPut state._write
    red = if count < state.red then 1 else 0
    green = if count < state.green then 1 else 0
    blue = if count < state.blue then 1 else 0

