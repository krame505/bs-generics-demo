package DemoSim where

import Demo
import UART
import RGB
import Buttons

import GetPut
import Connectable
import FIFO

{-# verilog sysDemoSim #-}
sysDemoSim :: Module Empty
sysDemoSim = module
  demo <- mkDemo

  tty <- mkReg InvalidFile
  init <- mkReg False

  rules
    "init": when not init ==> do
      fh <- $fopen "ttySim" "rb+"
      tty := fh
      init := True
    
    "tx": when True ==> do
      c <- demo.txData.get
      $display "Tx %x" c
      $fwrite tty "%c" (pack c)

    "rx": when True ==> do
      c <- $fgetc tty
      if c /= negate 1
        then do $display "Rx %x" c
                demo.rxData.put $ truncate $ pack c
        else noAction
