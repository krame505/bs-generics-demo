
import "BDPI" function ActionValue#(UInt#(32)) rxData();
import "BDPI" function Action txData(Bit#(8) data);
