-- Copyright 2021 Google LLC
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--      http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.

package UART where

import GetPut
import FIFOF

interface UART =
  txData :: Put (Bit 8)
  rxData :: Get (Bit 8)

  tx :: Bit 1
  rx :: Bit 1 -> Action

clockFreq :: Integer
clockFreq = 100000000

data State = Ready | StartBit | DataBit (UInt 3) | StopBit
  deriving (Eq, Bits)

mkUART :: Integer -> Module UART
mkUART baud = module
  let bitCounts = clockFreq / baud - 1
  let sampleCounts = bitCounts / 2

  txFIFO :: FIFOF (Bit 8) <- mkFIFOF
  txState :: Reg State <- mkReg Ready
  txCounter :: Reg (UInt 32) <- mkReg 0
  txBit :: Reg (Bit 1) <- mkReg 1

  rxFIFO :: FIFOF (Bit 8) <- mkFIFOF
  rxState :: Reg State <- mkReg Ready
  rxCounter :: Reg (UInt 32) <- mkReg 0
  rxByte :: Reg (Bit 8) <- mkReg 0
  rxBit :: Reg (Bit 1) <- mkReg 1

  rules
    "tx": when txCounter == 0 && txFIFO.notEmpty ==> do
      case txState of
        Ready -> do
          txState := StartBit
        StartBit -> do
          txState := DataBit 0
          txBit := 0
          txCounter := fromInteger bitCounts
        DataBit i -> do
          txState := if i == 7 then StopBit else DataBit (i + 1)
          txBit := truncate (txFIFO.first >> i)
          txCounter := fromInteger bitCounts
        StopBit -> do
          txState := Ready
          txBit := 1
          txFIFO.deq
          txCounter := fromInteger bitCounts

    "update_tx_counter": when txCounter > 0 ==>
      txCounter := txCounter - 1

    "rx": when rxCounter == 0 ==> do
      case rxState of
        Ready -> do
          rxState := StartBit
          rxCounter := fromInteger sampleCounts
        StartBit ->
          if rxBit == 0  -- Check start bit is 0
            then do
              rxState := DataBit 0
              rxCounter := fromInteger bitCounts
            else rxState := Ready
        DataBit i -> do
          rxState := if i == 7 then StopBit else DataBit (i + 1)
          rxByte := rxByte | (zeroExtend rxBit) << i
          rxCounter := fromInteger bitCounts
        StopBit -> do
          rxState := Ready
          if rxBit == 1  -- Check stop bit is 1
            then rxFIFO.enq rxByte
            else noAction
          rxByte := 0
          rxCounter := fromInteger sampleCounts

    "update_rx_counter": when rxCounter > 0 ==>
      rxCounter := rxCounter - 1

  interface
    txData = toPut txFIFO
    rxData = toGet rxFIFO
    tx = txBit
    rx = rxBit._write
