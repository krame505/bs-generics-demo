package SumSquares where

import CShow
import Vector
import FIFO
import GetPut

type Id = Bit 16 -- Try changing the size

-- Try adding/reordering constructors
data CounterCommand
  = Num (Int 32)
  | ResetSum
  | ResetSquareSum
  deriving (Bits)

struct CounterRequest =
  id :: Id
  command :: CounterCommand
 deriving (Bits)

struct CounterResponse a =
  id :: Id
  val :: a
 deriving (Bits)

interface Counter =
  requests :: Put CounterRequest
  sum :: Get (CounterResponse (Int 32))
  squareSum :: Get (CounterResponse (Int 64))

{-# verilog mkCounter #-}
mkCounter :: Module Counter
mkCounter = module
  requests <- mkFIFO
  sums <- mkFIFO
  squareSums <- mkFIFO

  sum :: Reg (Int 32) <- mkReg 0
  squareSum :: Reg (Int 64) <- mkReg 0

  rules
    "handle_request": when True ==> do
      -- $display "Handling request " (cshow requests.first)
      let newSum =
            case requests.first.command of
               Num n -> sum + n
               ResetSum -> 0
               _ -> sum
          newSquareSum =
            case requests.first.command of
               Num n -> squareSum + (signExtend n) * (signExtend n)
               ResetSquareSum -> 0
               _ -> squareSum
      sums.enq (CounterResponse { id = requests.first.id; val = newSum; })
      squareSums.enq (CounterResponse { id = requests.first.id; val = newSquareSum; })
      sum := newSum
      squareSum := newSquareSum
      requests.deq

  interface
    requests = toPut requests
    sum = toGet sums
    squareSum = toGet squareSums
