package Demo where

import GenCRepr
import GenCMsg
import CShow
import Vector
import GetPut
import Connectable
import UART
import COBS
import Counter
import RGB

type NumRGBs = 4

struct RGBCommand =
  addr :: UInt (TLog NumRGBs)
  state :: RGB
 deriving (Bits)

type NumButtons = 4

interface DemoMsgs =
  -- In order of highest to lowest urgency
  -- Try changing the order and FIFO sizes
  ctrCommands :: Rx 16 16 CounterCommand
  sums        :: Tx 16 2 (Result (Int 16))
  products    :: Tx 16 2 (Result (Int 64))

  rgbCommands :: Rx 8 8 RGBCommand

  buttonEvents :: Tx 8 8 (UInt NumButtons)

interface Top =
  tx :: Bit 1 {-# always_ready, always_enabled #-}
  rx :: Bit 1 -> Action {-# always_ready, always_enabled, prefix="", arg_names = [rx] #-}
  red :: Bit NumRGBs {-# always_ready, always_enabled #-}
  green :: Bit NumRGBs {-# always_ready, always_enabled #-}
  blue :: Bit NumRGBs {-# always_ready, always_enabled #-}
  buttons :: Bit NumButtons -> Action {-# always_ready, always_enabled, prefix="", arg_names = [buttons] #-}

{-# verilog mkTop #-}
mkTop :: Module Top
mkTop = mkTopReal

-- Seperated out due to the context...
mkTopReal :: (GenCMsg DemoMsgs rxBytes txBytes) => Module Top
mkTopReal = module
  writeCMsgDecls "demo" (_ :: DemoMsgs)

  uart <- mkUART 115200
  enc :: COBSEncoder txBytes <- mkCOBSEncoder
  dec :: COBSDecoder rxBytes <- mkCOBSDecoder
  msgMgr :: MsgManager DemoMsgs rxBytes txBytes <- mkMsgManager

  uart.rxData <-> dec.byte
  dec.msg <-> dropSize msgMgr.rxMsg
  msgMgr.txMsg <-> enc.msg
  enc.byte <-> uart.txData

  ctr <- mkCounter
  toGet msgMgr.fifos.ctrCommands <-> ctr.command
  ctr.sum <-> toPut msgMgr.fifos.sums
  ctr.product <-> toPut msgMgr.fifos.products

  rgbs :: Vector NumRGBs RGBControl <- replicateM mkRGBControl
  rules
    "write_rgb": when True ==> do
      let c = msgMgr.fifos.rgbCommands.first
      (select rgbs c.addr).state.put c.state
      msgMgr.fifos.rgbCommands.deq

  let buttonDebounce = 10000 -- Clock cycles to wait before declaring a press
  buttonCounts :: Vector NumButtons (Reg (UInt 16)) <- replicateM $ mkReg 0
  buttonSent :: Vector NumButtons (Reg Bool) <- replicateM $ mkReg False
  let readButtons :: Bit NumButtons -> Action
      readButtons x = mapM_
        (\ i ->
          if (1 & (x >> i)) == 1 && (buttonCounts !! i)._read <= maxBound
          then buttonCounts !! i := (buttonCounts !! i)._read + 1
          else do buttonCounts !! i := 0
                  buttonSent !! i := False
        )
        (genVector :: Vector NumButtons Integer)
  addRules $ foldr1 (<+) $ map
    (\ i ->
      rules
        ("send_button_" +++ integerToString i):
            when not (buttonSent !! i)._read && (buttonCounts !! i)._read >= buttonDebounce ==> do
          msgMgr.fifos.buttonEvents.enq (fromInteger i)
          buttonSent !! i := True
    )
    (genVector :: Vector NumButtons Integer)

  interface
    tx = uart.tx
    rx = uart.rx
    red = Prelude.pack $ map (\ c -> (c::RGBControl).red) rgbs
    green = Prelude.pack $ map (\ c -> (c::RGBControl).green) rgbs
    blue = Prelude.pack $ map (\ c -> (c::RGBControl).blue) rgbs
    buttons = readButtons
