package DemoSim where

import Demo
import PTY
import RGB
import Buttons

import GenCMsg
import COBS
import GetPut
import Connectable
import FIFO

interface DemoSimMsgs =
  rgbCommands :: Tx 8 8 (RGBCommand NumRGBs)
  buttonEvents :: Rx 8 8 (UInt (TLog NumButtons))

mkDemoSim :: (GenCMsg DemoSimMsgs rxBytes txBytes) => Module Empty
mkDemoSim = module
  writeCMsgDecls "demo_sim" (_ :: DemoSimMsgs)
  msgMgr :: MsgManager DemoSimMsgs rxBytes txBytes <- mkMsgManager
  enc :: COBSEncoder txBytes <- mkCOBSEncoder
  dec :: COBSDecoder rxBytes <- mkCOBSDecoder
  dec.msg <-> dropSize msgMgr.rxMsg
  msgMgr.txMsg <-> enc.msg

  demo <- mkDemo
  demo.rgbCommands <-> toPut msgMgr.fifos.rgbCommands
  toGet msgMgr.fifos.buttonEvents <-> demo.buttonEvents

  -- Wait for first byte to be recieved before sending data
  clientWriteEnable <- mkReg False
  simWriteEnable <- mkReg False

  rules
    "txClient": when clientWriteEnable ==> do
      c <- demo.txData.get
      -- $display "Tx %x" c
      txClient c

    "rxClient": when True ==> do
      c <- rxClient
      if c /= negate 1
        then do -- $display "Rx %x" ((truncate $ pack c) :: Bit 8)
                demo.rxData.put $ truncate $ pack c
                clientWriteEnable := True
        else noAction

    "txSim": when simWriteEnable ==> do
      c <- enc.byte.get
      txSim c

    "rxSim": when True ==> do
      c <- rxSim
      if c /= negate 1
        then do dec.byte.put $ truncate $ pack c
                simWriteEnable := True
        else noAction

{-# verilog sysDemoSim #-}
sysDemoSim :: Module Empty
sysDemoSim = mkDemoSim
